module length (
	input wire [31:0] op,
	output wire [5:0] op_length
);


assign op_length = (op[31:16] == 16'd0)? 
						(
							(op[15:8] == 8'd0)?
								(
									(op[7:4] == 4'd0)?
									(
										(op[3:2] == 2'd0)?
											(
												(op[1] == 1'd0)?op[0]:6'd2
											)
											:
											(
												(op[3] == 1'd0)?6'd3:6'd4
											)

									)
									:
									(
										(op[7:6] == 2'd0)?
											(
												(op[5] == 1'd0)?6'd5:6'd6
											)
											:
											(
												(op[7] == 1'd0)?6'd7:6'd8
											)
									)
								)
								:
								(
									(op[15:12] == 4'd0)?
									(
										(op[11:10] == 2'd0)?
											(
												(op[9] == 1'd0)?6'd9:6'd10
											)
											:
											(
												(op[11] == 1'd0)?6'd11:6'd12
											)

									)
									:
									(
										(op[15:14] == 2'd0)?
											(
												(op[13] == 1'd0)?6'd13:6'd14
											)
											:
											(
												(op[15] == 1'd0)?6'd15:6'd16
											)
									)
								) 
								
						)
						: 
						(
								(op[31:24] == 8'd0)?
								(
									(op[23:20] == 4'd0)?
									(
										(op[19:18] == 2'd0)?
											(
												(op[17] == 1'd0)?6'd17:6'd18
											)
											:
											(
												(op[19] == 1'd0)?6'd19:6'd20
											)

									)
									:
									(
										(op[23:22] == 2'd0)?
											(
												(op[21] == 1'd0)?6'd21:6'd22
											)
											:
											(
												(op[23] == 1'd0)?6'd23:6'd24
											)
									)
								)
								:
								(
									(op[31:28] == 4'd0)?
									(
										(op[27:26] == 2'd0)?
											(
												(op[25] == 1'd0)?6'd25:6'd26
											)
											:
											(
												(op[27] == 1'd0)?6'd27:6'd28
											)

									)
									:
									(
										(op[31:30] == 2'd0)?
											(
												(op[29] == 1'd0)?6'd29:6'd30
											)
											:
											(
												(op[31] == 1'd0)?6'd31:6'd32
											)
									)
								) 

						) ;

endmodule
