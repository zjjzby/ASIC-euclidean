module top(
		input wire [31:0] opa,
		input wire [31:0] opb,
		input wire start,
		input wire rst,
		input wire clk,
		output done,
		output [31:0] result
);

reg [2:0] current_state;
reg [2:0] next_state;
reg [31:0] regopa;
reg [31:0] regopb;

reg [31:0] result;
reg done;



reg [5:0] length_diff_reg;

wire [5:0] length_opa;
wire [5:0] length_opb;
wire [5:0] length_diff;

wire [31:0] length_in_opa;
wire [31:0] length_in_opb;
//***********************************************************************//
//                                                                       //
//                          state   machine                              //
//                                                                       //
//***********************************************************************//

parameter IDLE = 3'd0;
parameter INPUT = 3'd1;
parameter ADJUDICATE = 3'd2;
parameter CAMP_SWITCH = 3'd3;
parameter ALIGN = 3'd4;
parameter ABSOLUTE = 3'd5;
parameter OUTPUT = 3'd6;

parameter ZEROS = 32'd0;
parameter ZEROS_C = 7'b0; 


//***********************************************************************//
//                                                                       //
//                          state   machine                              //
//                                                                       //
//***********************************************************************//
always @(posedge clk or negedge rst) begin : proc_current_state
	if(~rst) begin
		current_state <= IDLE;
	end else begin
		current_state <= next_state ;
	end
end



always @ * begin : proc_next_state
	case (current_state)
		IDLE:begin 
			if(start == 1) 
				next_state <= INPUT;
			else 
				next_state <= IDLE;			
		end
		INPUT:next_state <= ADJUDICATE;
		ADJUDICATE:begin 
			if(regopa == regopb || regopa == 0 || regopb == 0) begin
				next_state <= OUTPUT;
			end
			else begin 
				next_state <= CAMP_SWITCH;
			end
		end
		CAMP_SWITCH:next_state <= ALIGN;
		ALIGN:next_state <= ABSOLUTE;
		ABSOLUTE:next_state <= ADJUDICATE;
		OUTPUT:begin 
			if(start == 1) 
				next_state <= INPUT;
			else 
				next_state <= IDLE;
		end
		default : next_state <= IDLE;
	endcase
end



//***********************************************************************//
//                                                                       //
//                                                                       //
//                                                                       //
//***********************************************************************//
always @(posedge clk or negedge rst) begin : proc_regopa
	if(~rst) begin
		regopa <= ZEROS;
	end else begin
		case (next_state)
			IDLE:regopa <= ZEROS;
			INPUT:regopa <= opa;
			ADJUDICATE:regopa <= regopa;
			CAMP_SWITCH:begin 
				if(regopa < regopb) begin
					regopa <= regopb;
				end
				else begin 
					regopa <= regopa;
				end
			end
			ALIGN:regopa <= regopa;
			ABSOLUTE:begin 
				if (regopa >= regopb ) begin 
					regopa <= regopa - regopb;
				end
				else begin 
					regopa <= regopb - regopa;
				end
			end		
			default :regopa <= regopa;
		endcase		
	end
end

//

always @(posedge clk or negedge rst) begin : proc_regopb
	if(~rst) begin
		regopb <= ZEROS;
	end else begin
		case (next_state)
			IDLE:regopb <= ZEROS;
			INPUT:regopb <= opb;
			ADJUDICATE:regopb <= regopb;
			CAMP_SWITCH:begin 
				if(regopa < regopb) begin
					regopb <= regopa <<< length_diff;
				end
				else begin 
					regopb <= regopb <<< length_diff;
				end
			end
			ALIGN:regopb <= regopb ;
			ABSOLUTE:regopb <= regopb >>> length_diff_reg;
			default:regopb <= regopb;
		endcase		
	end
end






assign length_in_opa = regopa;
assign length_in_opb = regopb;

length cal_opa_length(.op(length_in_opa), .op_length(length_opa));
length cal_opp_length(.op(length_in_opb), .op_length(length_opb));

assign length_diff = (length_opa >= length_opb)? (length_opa - length_opb):(length_opb - length_opa);



always @(posedge clk or negedge rst) begin : proc_length_diff_reg
	if(~rst) begin
		length_diff_reg <= 0;
	end else begin
		case (next_state)
			CAMP_SWITCH:begin 
				length_diff_reg <= length_diff;
			end
			default : length_diff_reg <= length_diff_reg;
		endcase
	end
end






//***********************************************************************//
//                                                                       //
//                       result                                          //
//                                                                       //
//***********************************************************************//


always @(posedge clk or negedge rst) begin : proc_result
	if(~rst) begin
		result <= ZEROS;
	end else begin
		case (next_state)
			OUTPUT:begin 
				if(regopa == regopb) begin 
					result <= regopa ;
				end
				else if (regopa == 0 ) begin
					result <=  regopb ;
				end
				else begin 
					result <= regopa ;
				end
			end
			default : begin 
				result <= result;
			end
		endcase
	end
end


always @(posedge clk or negedge rst) begin : proc_done
	if(~rst) begin
		done <= 1'b0;
	end else begin
		case (next_state)
			OUTPUT: begin 
				done <= 1'b1;
			end
			default : done <= 1'b0;
		endcase
	end
end


endmodule // top
